
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Calculates the ppb error from expected count.
-- 
-- Input is count in the expected frequency g_frequency over one second.
-- The measurement period 1s is expected to be correct.
entity freq_offset_from_count is
    generic (
        g_frequency : in real
    );
    port (
        clk_i: in std_logic;
        count_i: in unsigned(31 downto 0);
        count_vld_i: in std_logic;
        error_ppb_o : out integer range -10000 to 10000;
        error_ppb_vld_o : out std_logic
        );
end freq_offset_from_count;

architecture rtl of freq_offset_from_count is

    constant c_expected_count : unsigned(31 downto 0) := to_unsigned(natural(g_frequency), 32);
    constant c_ppm : integer range 0 to 100 := natural(g_frequency/1.0e6);
    
    signal offset : integer range -10000 to 10000 := 0;
    signal error_ppb : integer range -10000 to 10000 := 0;

    type state_type is (idle, calc_error, output_error);
    signal state : state_type := idle;
begin

    p_error : process (clk_i)
    begin
        if rising_edge(clk_i) then
            error_ppb_vld_o <= '0';
            case state is
                when idle =>
                    if count_vld_i = '1' then
                        state <= calc_error;
                        offset <= to_integer(count_i - c_expected_count);
                    end if;

                when calc_error =>
                    state <= output_error;
                    error_ppb <= offset * 1000 / c_ppm;

                when output_error =>
                    state <= idle;
                    error_ppb_o <= error_ppb;
                    error_ppb_vld_o <= '1';
            end case;
        end if;
    end process;
    

end rtl;