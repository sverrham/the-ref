
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity freq_offset_from_count is
    generic (
        g_frequency : in real
    );
    port (
        i_clk: in std_logic;
        i_count: in unsigned(31 downto 0);
        i_count_vld: in std_logic;
        o_error_ppm : out integer range -255 to 256;
        o_error_ppm_vld : out std_logic
        );
end freq_offset_from_count;

architecture rtl of freq_offset_from_count is

    constant c_expected_count : unsigned(31 downto 0) := to_unsigned(natural(g_frequency), 32);
    constant c_ppm : integer range 0 to 100 := natural(g_frequency/1.0e6);
    
    signal offset : integer range -1023 to 1024 := 0;
    signal error_ppm : integer range -1023 to 1024 := 0;

    type state_type is (idle, calc_error, output_error);
    signal state : state_type := idle;
begin

    p_error : process (i_clk)
    begin
        if rising_edge(i_clk) then
            o_error_ppm_vld <= '0';
            case state is
                when idle =>
                    if i_count_vld = '1' then
                        state <= calc_error;
                        offset <= to_integer(i_count - c_expected_count);
                    end if;

                when calc_error =>
                    state <= output_error;
                    error_ppm <= offset / c_ppm;

                when output_error =>
                    state <= idle;
                    o_error_ppm <= error_ppm;
                    o_error_ppm_vld <= '1';
            end case;
        end if;
    end process;
    

end rtl;